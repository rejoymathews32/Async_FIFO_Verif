// Author - Rejoy Roy Mathews
// Modify the parameter definitions in this file to test different Asynchronous
// FIFO configurations

localparam FIFO_DATA_WIDTH = 32;
localparam FIFO_DEPTH = 8;
localparam SYNCHRONIZER_FLOPS = 2;
